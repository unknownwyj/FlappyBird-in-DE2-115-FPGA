module decodecolor(input [7:0]color, output [7:0]red, output [7:0]green, output [7:0]blue);
    wire [23:0]colormap[0:255];
    assign colormap[0] = 24'h543847;
    assign colormap[1] = 24'h000000;
    assign colormap[2] = 24'h533846;
    assign colormap[3] = 24'h54d1ff;
    assign colormap[4] = 24'hfafafa;
    assign colormap[5] = 24'h4bc1f8;
    assign colormap[6] = 24'hd7e6cc;
    assign colormap[7] = 24'hfcd884;
    assign colormap[8] = 24'he46018;
    assign colormap[9] = 24'h40a4d2;
    assign colormap[10] = 24'hffffff;
    assign colormap[11] = 24'he4fd8b;
    assign colormap[12] = 24'h73bf2e;
    assign colormap[13] = 24'h9ce659;
    assign colormap[14] = 24'h558022;
    assign colormap[15] = 24'hd7a84c;
    assign colormap[16] = 24'hded895;
    assign colormap[17] = 24'hffffff;
    assign colormap[18] = 24'h000000;
    assign colormap[19] = 24'h533846;
    assign colormap[20] = 24'hfc730f;
    assign colormap[21] = 24'hfafafa;
    assign colormap[22] = 24'hfc3800;
    assign colormap[23] = 24'hd7e6cc;
    assign colormap[24] = 24'hf8b733;
    assign colormap[25] = 24'hd32f00;
    assign colormap[26] = 24'hffffff;
    assign colormap[27] = 24'h543847;
    assign colormap[28] = 24'h523745;
    assign colormap[29] = 24'h00a848;
    assign colormap[30] = 24'h58d858;
    assign colormap[31] = 24'hff290d;
    assign colormap[32] = 24'hffffff;
    assign colormap[33] = 24'hfafafa;
    assign colormap[34] = 24'hd6d6d6;
    assign colormap[35] = 24'hffffff;
    assign colormap[36] = 24'h000000;
    assign colormap[37] = 24'hfc730f;
    assign colormap[38] = 24'hfafafa;
    assign colormap[39] = 24'hfc3800;
    assign colormap[40] = 24'hd7e6cc;
    assign colormap[41] = 24'hf8b733;
    assign colormap[42] = 24'hd32f00;
    assign colormap[43] = 24'hffffff;
    assign colormap[44] = 24'h008793;
    assign colormap[45] = 24'haee8d2;
    assign colormap[46] = 24'h00b3c2;
    assign colormap[47] = 24'h00818c;
    assign colormap[48] = 24'h0093a0;
    assign colormap[49] = 24'hfcb800;
    assign colormap[50] = 24'h00b200;
    assign colormap[51] = 24'h00a300;
    assign colormap[52] = 24'hffffff;
    assign colormap[53] = 24'hffffff;
    assign colormap[54] = 24'h543847;
    assign colormap[55] = 24'hc0dd71;
    assign colormap[56] = 24'hd9f383;
    assign colormap[57] = 24'he4fd8b;
    assign colormap[58] = 24'hdff987;
    assign colormap[59] = 24'haccc62;
    assign colormap[60] = 24'ha2c35a;
    assign colormap[61] = 24'h8db14b;
    assign colormap[62] = 24'h799f3d;
    assign colormap[63] = 24'h709836;
    assign colormap[64] = 24'h608a2a;
    assign colormap[65] = 24'h5a8426;
    assign colormap[66] = 24'h558022;
    assign colormap[67] = 24'hd1ed7d;
    assign colormap[68] = 24'hdff988;
    assign colormap[69] = 24'hd9f483;
    assign colormap[70] = 24'hc9e577;
    assign colormap[71] = 24'h79a03c;
    assign colormap[72] = 24'h67912f;
    assign colormap[73] = 24'hd1ec7d;
    assign colormap[74] = 24'hc9e678;
    assign colormap[75] = 24'h98ba52;
    assign colormap[76] = 24'h709736;
    assign colormap[77] = 24'hc4e173;
    assign colormap[78] = 24'hdcf685;
    assign colormap[79] = 24'hb5d368;
    assign colormap[80] = 24'h689130;
    assign colormap[81] = 24'h5d8728;
    assign colormap[82] = 24'hb5d468;
    assign colormap[83] = 24'hd0ec7d;
    assign colormap[84] = 24'hc3e073;
    assign colormap[85] = 24'ha4c55c;
    assign colormap[86] = 24'h94b851;
    assign colormap[87] = 24'h84a945;
    assign colormap[88] = 24'h769c3a;
    assign colormap[89] = 24'h000000;
    assign colormap[90] = 24'h533846;
    assign colormap[91] = 24'hfad78c;
    assign colormap[92] = 24'hfafafa;
    assign colormap[93] = 24'hf8b733;
    assign colormap[94] = 24'hd7e6cc;
    assign colormap[95] = 24'hfc3800;
    assign colormap[96] = 24'he0802c;
    assign colormap[97] = 24'hffffff;
    assign colormap[98] = 24'h94b751;
    assign colormap[99] = 24'ha5c65c;
    assign colormap[100] = 24'hdbf685;
    assign colormap[101] = 24'hc4e174;
    assign colormap[102] = 24'h5d8828;
    assign colormap[103] = 24'hc3e074;
    assign colormap[104] = 24'h000000;
    assign colormap[105] = 24'h533846;
    assign colormap[106] = 24'hfad78c;
    assign colormap[107] = 24'hfafafa;
    assign colormap[108] = 24'hf8b733;
    assign colormap[109] = 24'hd7e6cc;
    assign colormap[110] = 24'hfc3800;
    assign colormap[111] = 24'he0802c;
    assign colormap[112] = 24'hffffff;
    assign colormap[113] = 24'h000000;
    assign colormap[114] = 24'h533846;
    assign colormap[115] = 24'hfc730f;
    assign colormap[116] = 24'hfafafa;
    assign colormap[117] = 24'hfc3800;
    assign colormap[118] = 24'hd7e6cc;
    assign colormap[119] = 24'hf8b733;
    assign colormap[120] = 24'hd32f00;
    assign colormap[121] = 24'hffffff;
    assign colormap[122] = 24'hb8e6c4;
    assign colormap[123] = 24'he1f9d8;
    assign colormap[124] = 24'h54c4cc;
    assign colormap[125] = 24'h9ddbd5;
    assign colormap[126] = 24'hd9f6d7;
    assign colormap[127] = 24'hd2efc6;
    assign colormap[128] = 24'h97d9d3;
    assign colormap[129] = 24'hcdecc4;
    assign colormap[130] = 24'h5ce16f;
    assign colormap[131] = 24'h65c9cc;
    assign colormap[132] = 24'ha1dcd7;
    assign colormap[133] = 24'hade4bd;
    assign colormap[134] = 24'hddefcf;
    assign colormap[135] = 24'hc5ebbc;
    assign colormap[136] = 24'hd0edc8;
    assign colormap[137] = 24'h5dcb79;
    assign colormap[138] = 24'hdaedce;
    assign colormap[139] = 24'h5adf6f;
    assign colormap[140] = 24'hd5f0c6;
    assign colormap[141] = 24'he7fbd9;
    assign colormap[142] = 24'h52cb6c;
    assign colormap[143] = 24'h67cc7f;
    assign colormap[144] = 24'h62df75;
    assign colormap[145] = 24'he1f1d0;
    assign colormap[146] = 24'he5fad8;
    assign colormap[147] = 24'he9fcd9;
    assign colormap[148] = 24'h5ee270;
    assign colormap[149] = 24'h4ec0ca;
    assign colormap[150] = 24'hffa791;
    assign colormap[151] = 24'he08b6b;
    assign colormap[152] = 24'hd78363;
    assign colormap[153] = 24'hbe744f;
    assign colormap[154] = 24'hb66f48;
    assign colormap[155] = 24'h8f5629;
    assign colormap[156] = 24'hfe9d82;
    assign colormap[157] = 24'hf09377;
    assign colormap[158] = 24'hf6987d;
    assign colormap[159] = 24'h9e5f36;
    assign colormap[160] = 24'hffa189;
    assign colormap[161] = 24'hc57a55;
    assign colormap[162] = 24'hec9173;
    assign colormap[163] = 24'hffa085;
    assign colormap[164] = 24'hec9273;
    assign colormap[165] = 24'hde8869;
    assign colormap[166] = 24'hac6a3f;
    assign colormap[167] = 24'h9f6136;
    assign colormap[168] = 24'h965a2e;
    assign colormap[169] = 24'hb76f49;
    assign colormap[170] = 24'hc47754;
    assign colormap[171] = 24'hd17f5e;
    assign colormap[172] = 24'hdf8a69;
    assign colormap[173] = 24'hab673f;
    assign colormap[174] = 24'hb87049;
    assign colormap[175] = 24'hd2815e;
    assign colormap[176] = 24'heb9073;
    assign colormap[177] = 24'hde8a6a;
    assign colormap[178] = 24'hea9174;
    assign colormap[179] = 24'hFFFFFF; // white 
    assign colormap[180] = 24'hf0e9a5;
    assign colormap[181] = 24'hc7c189;
    assign colormap[182] = 24'he8a147;
    assign colormap[183] = 24'he9e1e1;
    assign colormap[184] = 24'h9e9898;
    assign colormap[185] = 24'hc8c0c0;
    assign colormap[186] = 24'h847f7f;
    assign colormap[187] = 24'hedf16b;
    assign colormap[188] = 24'hbda14e;
    assign colormap[189] = 24'hfeda68;
    assign colormap[190] = 24'he2c25e;
    assign colormap[191] = 24'hf9f7f7;
    assign colormap[192] = 24'hd0cece;
    assign colormap[193] = 24'h878686;
    assign colormap[194] = 24'hefeded;
    assign colormap[195] = 24'hdf7126;// flame
    assign colormap[196] = 24'hfbf236;// flame
    assign colormap[254] = 24'hFFFFFF;
	assign colormap[255] = 24'hFFFFFF;
    assign {red, green, blue} = colormap[color];
endmodule